module tvxml

