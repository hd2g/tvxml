module xml

fn test_dummy() {
  assert true
}
